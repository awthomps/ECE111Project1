module fibonacci_calculator(input_s, reset_n, begin_fibo, clk, done, fibo_out);
	input [4:0] input_s;
	input reset_n;
	input begin_fibo; //Start calculation
	input clk;
	
	output done;
	output [15:0] fibo_out;
	
	


endmodule